module INSTR // a synthesisable rom implementation
(
	input [31:0] pc,
	output [31:0] instruction
);
	/* lw $3, 0($0) --
	Loop: slti $1, $3, 50
	beq $1, $0, Skip
	add $4, $4, $3
	addi $3, $3, 1
	beq $0, $0, Loop--
	Skip
	*/
	wire [29:0] i = pc[31:2];
	reg [31:0] rom[16:1];
	initial
	begin
		rom[1] = 32'b101000_10001_10001_0000000000010001; // #addi $s1, $s1, 17 PC 4
		rom[2] = 32'b101000_00011_00011_0000000000000011; // #addi $s2, $s2, 3 PC 8
		rom[3] = 32'b101000_00011_01000_00000_00000_000000; // #addi $t1, $s2, 0 PC 12
		rom[4] = 32'b000000_10001_01000_01001_00000_100010; // #sub $t2, $s1, $t1 PC 16
		rom[5] = 32'b000000_10001_01000_01010_00000_101010; // #slt $t3, $s1, $t1 PC 20
		rom[6] = 32'b000100_10001_01000_0000000000000100; // #beq $s1, $t1, 4 PC 24
		rom[7] = 32'b000110_01010_01011_0000000000000010; // #bne $t4, $t3, 2 PC 28
		rom[8] = 32'b000000_01000_00011_01000_00000_100000; // #add $t1, $t1, $s2 PC 32
		rom[9] = 32'b100110_00000000000000000000000100; // #jump 4 PC 36
		rom[10] = 32'b000000_01001_00011_01001_00000_100000; // #add $t2, $t2, $s2 PC 40
		rom[11] = 32'b101011_00011_01001_00000_00000_001000; // #sw $t2, 8($s2) PC 44
	end
	assign instruction = (pc < 48 )? rom[i]: 32'd0;
endmodule